library verilog;
use verilog.vl_types.all;
entity DM_tb is
end DM_tb;
