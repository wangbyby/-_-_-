library verilog;
use verilog.vl_types.all;
entity GPR_tb is
end GPR_tb;
