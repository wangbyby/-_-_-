library verilog;
use verilog.vl_types.all;
entity Controll_tb is
end Controll_tb;
