library verilog;
use verilog.vl_types.all;
entity MUX is
    port(
        a               : in     vl_logic_vector(31 downto 0);
        b               : in     vl_logic_vector(31 downto 0);
        choose          : in     vl_logic;
        z               : out    vl_logic_vector(31 downto 0)
    );
end MUX;
